

package test_lib_pkg;

  import uvm_pkg::*;
	
  `include "uvm_macros.svh"
  `include "axi_transaction.sv"
  `include "apb_transaction.sv"
  `include "axi_sequencer.sv"
  `include "axi_sequence.sv"
  `include "axi_monitor.sv"
  `include "apb_monitor.sv"
  `include "axi_driver.sv"
  `include "scoreboard.sv"
  `include "axi_agent.sv"
  `include "apb_agent.sv"
  `include "axi2apb_env.sv"
  `include "axi2apb_base_test.sv"


endpackage 
